// 
// Copyright 2020 Datum Technology Corporation
// 
// Licensed under the Solderpad Hardware License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     https://solderpad.org/licenses/
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 


`ifndef __UVMA_AXIS_MACROS_SV__
`define __UVMA_AXIS_MACROS_SV__


`define UVMA_AXIS_TDATA_MAX_SIZE  1_024
`define UVMA_AXIS_TID_MAX_SIZE        8
`define UVMA_AXIS_TDEST_MAX_SIZE      4
`define UVMA_AXIS_TUSER_MAX_SIZE  1_024


`endif // __UVMA_AXIS_MACROS_SV__
