// 
// Copyright 2020 Datum Technology Corporation
// 
// Licensed under the Solderpad Hardware License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     https://solderpad.org/licenses/
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 


`ifndef __UVMA_AXIS_MSTR_BASE_SEQ_SV__
`define __UVMA_AXIS_MSTR_BASE_SEQ_SV__


/**
 * TODO Describe uvma_axis_mstr_base_seq_c
 */
class uvma_axis_mstr_base_seq_c extends uvma_axis_base_seq_c;
   
   `uvm_object_utils(uvma_axis_mstr_base_seq_c)
   
   
   /**
    * Default constructor.
    */
   extern function new(string name="uvma_axis_mstr_base_seq");
   
endclass : uvma_axis_mstr_base_seq_c


function uvma_axis_mstr_base_seq_c::new(string name="uvma_axis_mstr_base_seq");
   
   super.new(name);
   
endfunction : new


`endif // __UVMA_AXIS_MSTR_BASE_SEQ_SV__
